library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Lab_2 is
port(a, b : in std_logic;
		f: out std_logic);
end Lab_2;

architecture Lab_2_arc of Lab_2 is
begin
		
end Lab_2_arc;